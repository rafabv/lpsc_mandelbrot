//--------------------------------------------------------------------------------
//                                 _             _
//                                | |_  ___ _ __(_)__ _
//                                | ' \/ -_) '_ \ / _` |
//                                |_||_\___| .__/_\__,_|
//                                         |_|
//
//--------------------------------------------------------------------------------
//
// Company: hepia
// Author: <author>
//
// Module Name: <prj_name>
// Target Device: <board_name> <part_name>
// Tool version: <tool_version>
// Description: <prj_name>
//
// Last update: <update_time>
//
//-------------------------------------------------------------------------------

package <prj_name>;
    
endpackage
