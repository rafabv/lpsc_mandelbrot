----------------------------------------------------------------------------------
--                                 _             _
--                                | |_  ___ _ __(_)__ _
--                                | ' \/ -_) '_ \ / _` |
--                                |_||_\___| .__/_\__,_|
--                                         |_|
--
----------------------------------------------------------------------------------
--
-- Company: hepia
-- Author: Joachim Schmidt <joachim.schmidt@hesge.ch>
--
-- Module Name: tb_lpsc_hdmi_interface_pkg - arch
-- Target Device:  xc7a200tsbg484-1
-- Tool version: 2021.2
-- Description: Testbench for package lpsc_hdmi_interface_pkg
--
-- Last update: 2022-02-28 08:45:30
--
---------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tb_lpsc_hdmi_interface_pkg is
end tb_lpsc_hdmi_interface_pkg;


architecture behavioral of tb_lpsc_hdmi_interface_pkg is

begin

end behavioral;
