----------------------------------------------------------------------------------
--                                 _             _
--                                | |_  ___ _ __(_)__ _
--                                | ' \/ -_) '_ \ / _` |
--                                |_||_\___| .__/_\__,_|
--                                         |_|
--
----------------------------------------------------------------------------------
--
-- Company: hepia
-- Author: <author>
--
-- Module Name: tb_<prj_name> - arch
-- Target Device: <board_name> <part_name>
-- Tool version: <tool_version>
-- Description: Testbench for package <prj_name>
--
-- Last update: <update_time>
--
---------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tb_<prj_name> is
end tb_<prj_name>;


architecture behavioral of tb_<prj_name> is

begin

end behavioral;
