----------------------------------------------------------------------------------
--                                 _             _
--                                | |_  ___ _ __(_)__ _
--                                | ' \/ -_) '_ \ / _` |
--                                |_||_\___| .__/_\__,_|
--                                         |_|
--
----------------------------------------------------------------------------------
--
-- Company: hepia
-- Author: <author>
--
-- Module Name: <prj_name> - arch
-- Target Device: <board_name> <part_name>
-- Tool version: <tool_version>
-- Description: Package <prj_name>
--
-- Last update: <update_time>
--
---------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package <prj_name> is

end <prj_name>;


package body <prj_name> is

end <prj_name>;
