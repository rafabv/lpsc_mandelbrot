//--------------------------------------------------------------------------------
//                                 _             _
//                                | |_  ___ _ __(_)__ _
//                                | ' \/ -_) '_ \ / _` |
//                                |_||_\___| .__/_\__,_|
//                                         |_|
//
//--------------------------------------------------------------------------------
//
// Company: hepia
// Author: <author>
//
// Module Name: tb_<prj_name> - arch
// Target Device: <board_name> <part_name>
// Tool version: <tool_version>
// Description: Testbench for <prj_name>
//
// Last update: <update_time>
//
//-------------------------------------------------------------------------------
`timescale 1ns / 1ps

import <prj_name>::*;

module tb_<prj_name> ();

// Stimulis generator
initial begin
  $finish;
end

endmodule
